`timescale 1ns / 1ps
module Instruction_Memory(
    input [63:0]Instr_Address,
    input reset,
    input clk, IF_ID_write,
    output reg [31:0]Instruction
    );
    reg[7:0]Ins_Reg[263:0];
    initial begin
Ins_Reg[0] = 8'h01;
Ins_Reg[1] = 8'h40; 
Ins_Reg[2] = 8'h05; 
Ins_Reg[3] = 8'h13; 
Ins_Reg[4] = 8'h00; 
Ins_Reg[5] = 8'h00; 
Ins_Reg[6] = 8'h04; 
Ins_Reg[7] = 8'h13; 
Ins_Reg[8] = 8'h00; 
Ins_Reg[9] = 8'h40; 
Ins_Reg[10] = 8'h05;
Ins_Reg[11] = 8'h93;
Ins_Reg[12] = 8'h00;
Ins_Reg[13] = 8'h50;
Ins_Reg[14] = 8'h02;
Ins_Reg[15] = 8'h93;
Ins_Reg[16] = 8'h00;
Ins_Reg[17] = 8'h40;
Ins_Reg[18] = 8'h0f;
Ins_Reg[19] = 8'h13;
Ins_Reg[20] = 8'h00;
Ins_Reg[21] = 8'h30;
Ins_Reg[22] = 8'h03;
Ins_Reg[23] = 8'h13;
Ins_Reg[24] = 8'h00;
Ins_Reg[25] = 8'h20;
Ins_Reg[26] = 8'h03;
Ins_Reg[27] = 8'h93;
Ins_Reg[28] = 8'h00;
Ins_Reg[29] = 8'h55;
Ins_Reg[30] = 8'h20;
Ins_Reg[31] = 8'h23;
Ins_Reg[32] = 8'h01;
Ins_Reg[33] = 8'he5;
Ins_Reg[34] = 8'h24;
Ins_Reg[35] = 8'h23;
Ins_Reg[36] = 8'h00;
Ins_Reg[37] = 8'h65;
Ins_Reg[38] = 8'h28;
Ins_Reg[39] = 8'h23;
Ins_Reg[40] = 8'h00;
Ins_Reg[41] = 8'h75;
Ins_Reg[42] = 8'h2c;
Ins_Reg[43] = 8'h23;
Ins_Reg[44] = 8'h00;
Ins_Reg[45] = 8'h00;
Ins_Reg[46] = 8'h80;
Ins_Reg[47] = 8'h93;
Ins_Reg[48] = 8'h00;
Ins_Reg[49] = 8'h00;
Ins_Reg[50] = 8'h80;
Ins_Reg[51] = 8'h93;
Ins_Reg[52] = 8'h00;
Ins_Reg[53] = 8'h00;
Ins_Reg[54] = 8'h80;
Ins_Reg[55] = 8'h93;
Ins_Reg[56] = 8'h00;
Ins_Reg[57] = 8'h04;
Ins_Reg[58] = 8'h0f;
Ins_Reg[59] = 8'h13;
Ins_Reg[60] = 8'h00;
Ins_Reg[61] = 8'h34;
Ins_Reg[62] = 8'h1e;
Ins_Reg[63] = 8'h93;
Ins_Reg[64] = 8'h00;
Ins_Reg[65] = 8'hae;
Ins_Reg[66] = 8'h8e;
Ins_Reg[67] = 8'hb3;
Ins_Reg[68] = 8'h08;
Ins_Reg[69] = 8'hb4;
Ins_Reg[70] = 8'h0e;
Ins_Reg[71] = 8'h63;
Ins_Reg[72] = 8'h00;
Ins_Reg[73] = 8'h00;
Ins_Reg[74] = 8'h80;
Ins_Reg[75] = 8'h93;
Ins_Reg[76] = 8'h00;
Ins_Reg[77] = 8'h00;
Ins_Reg[78] = 8'h80;
Ins_Reg[79] = 8'h93;
Ins_Reg[80] = 8'h00;
Ins_Reg[81] = 8'h00;
Ins_Reg[82] = 8'h80;
Ins_Reg[83] = 8'h93;
Ins_Reg[84] = 8'h00;
Ins_Reg[85] = 8'h00;
Ins_Reg[86] = 8'h80;
Ins_Reg[87] = 8'h93;
Ins_Reg[88] = 8'h00;
Ins_Reg[89] = 8'h00;
Ins_Reg[90] = 8'h80;
Ins_Reg[91] = 8'h93;
Ins_Reg[92] = 8'h00;
Ins_Reg[93] = 8'h00;
Ins_Reg[94] = 8'h80;
Ins_Reg[95] = 8'h93;
Ins_Reg[96] = 8'h00;
Ins_Reg[97] = 8'h3f;
Ins_Reg[98] = 8'h13;
Ins_Reg[99] = 8'h13;
Ins_Reg[100] = 8'h00;
Ins_Reg[101] = 8'h65;
Ins_Reg[102] = 8'h03;
Ins_Reg[103] = 8'h33;
Ins_Reg[104] = 8'h00;
Ins_Reg[105] = 8'h0e;
Ins_Reg[106] = 8'ha3;
Ins_Reg[107] = 8'h83;
Ins_Reg[108] = 8'h00;
Ins_Reg[109] = 8'h0f;
Ins_Reg[110] = 8'h8f;
Ins_Reg[111] = 8'h93;
Ins_Reg[112] = 8'h00;
Ins_Reg[113] = 8'h03;
Ins_Reg[114] = 8'h2e;
Ins_Reg[115] = 8'h03;
Ins_Reg[116] = 8'h00;
Ins_Reg[117] = 8'h0f;
Ins_Reg[118] = 8'h8f;
Ins_Reg[119] = 8'h93;
Ins_Reg[120] = 8'h04;
Ins_Reg[121] = 8'h7e;
Ins_Reg[122] = 8'h42;
Ins_Reg[123] = 8'h63;
Ins_Reg[124] = 8'h00;
Ins_Reg[125] = 8'h00;
Ins_Reg[126] = 8'h80;
Ins_Reg[127] = 8'h93;
Ins_Reg[128] = 8'h00;
Ins_Reg[129] = 8'h00;
Ins_Reg[130] = 8'h80;
Ins_Reg[131] = 8'h93;
Ins_Reg[132] = 8'h00;
Ins_Reg[133] = 8'h00;
Ins_Reg[134] = 8'h80;
Ins_Reg[135] = 8'h93;
Ins_Reg[136] = 8'h00;
Ins_Reg[137] = 8'h00;
Ins_Reg[138] = 8'h80;
Ins_Reg[139] = 8'h93;
Ins_Reg[140] = 8'h00;
Ins_Reg[141] = 8'h00;
Ins_Reg[142] = 8'h80;
Ins_Reg[143] = 8'h93;
Ins_Reg[144] = 8'h00;
Ins_Reg[145] = 8'h00;
Ins_Reg[146] = 8'h80;
Ins_Reg[147] = 8'h93;
Ins_Reg[148] = 8'h00;
Ins_Reg[149] = 8'h1f;
Ins_Reg[150] = 8'h0f;
Ins_Reg[151] = 8'h13;
Ins_Reg[152] = 8'hfa;
Ins_Reg[153] = 8'hbf;
Ins_Reg[154] = 8'h4e;
Ins_Reg[155] = 8'he3;
Ins_Reg[156] = 8'h00;
Ins_Reg[157] = 8'h00;
Ins_Reg[158] = 8'h80;
Ins_Reg[159] = 8'h93;
Ins_Reg[160] = 8'h00;
Ins_Reg[161] = 8'h00;
Ins_Reg[162] = 8'h80;
Ins_Reg[163] = 8'h93;
Ins_Reg[164] = 8'h00;
Ins_Reg[165] = 8'h00;
Ins_Reg[166] = 8'h80;
Ins_Reg[167] = 8'h93;
Ins_Reg[168] = 8'h00;
Ins_Reg[169] = 8'h14;
Ins_Reg[170] = 8'h04;
Ins_Reg[171] = 8'h13;
Ins_Reg[172] = 8'hf8;
Ins_Reg[173] = 8'h00;
Ins_Reg[174] = 8'h00;
Ins_Reg[175] = 8'he3;
Ins_Reg[176] = 8'h00;
Ins_Reg[177] = 8'h00;
Ins_Reg[178] = 8'h80;
Ins_Reg[179] = 8'h93;
Ins_Reg[180] = 8'h00;
Ins_Reg[181] = 8'h00;
Ins_Reg[182] = 8'h80;
Ins_Reg[183] = 8'h93;
Ins_Reg[184] = 8'h00;
Ins_Reg[185] = 8'h00;
Ins_Reg[186] = 8'h80;
Ins_Reg[187] = 8'h93;
Ins_Reg[188] = 8'h00;
Ins_Reg[189] = 8'h00;
Ins_Reg[190] = 8'h80;
Ins_Reg[191] = 8'h93;
Ins_Reg[192] = 8'h00;
Ins_Reg[193] = 8'h00;
Ins_Reg[194] = 8'h80;
Ins_Reg[195] = 8'h93;
Ins_Reg[196] = 8'h00;
Ins_Reg[197] = 8'h00;
Ins_Reg[198] = 8'h80;
Ins_Reg[199] = 8'h93;
Ins_Reg[200] = 8'h00;
Ins_Reg[201] = 8'h73;
Ins_Reg[202] = 8'h20;
Ins_Reg[203] = 8'h23;
Ins_Reg[204] = 8'h01;
Ins_Reg[205] = 8'hce;
Ins_Reg[206] = 8'ha0;
Ins_Reg[207] = 8'h23;
Ins_Reg[208] = 8'hfa;
Ins_Reg[209] = 8'h00;
Ins_Reg[210] = 8'h0c;
Ins_Reg[211] = 8'he3;
Ins_Reg[212] = 8'h00;
Ins_Reg[213] = 8'h00;
Ins_Reg[214] = 8'h80;
Ins_Reg[215] = 8'h93;
Ins_Reg[216] = 8'h00;
Ins_Reg[217] = 8'h00;
Ins_Reg[218] = 8'h80;
Ins_Reg[219] = 8'h93;
Ins_Reg[220] = 8'h00;
Ins_Reg[221] = 8'h00;
Ins_Reg[222] = 8'h80;
Ins_Reg[223] = 8'h93;
Ins_Reg[224] = 8'h00;
Ins_Reg[225] = 8'h00;
Ins_Reg[226] = 8'h80;
Ins_Reg[227] = 8'h93;
Ins_Reg[228] = 8'h00;
Ins_Reg[229] = 8'h00;
Ins_Reg[230] = 8'h80;
Ins_Reg[231] = 8'h93;
Ins_Reg[232] = 8'h00;
Ins_Reg[233] = 8'h00;
Ins_Reg[234] = 8'h80;
Ins_Reg[235] = 8'h93;
Ins_Reg[236] = 8'h00;
Ins_Reg[237] = 8'h05;
Ins_Reg[238] = 8'h22;
Ins_Reg[239] = 8'h83;
Ins_Reg[240] = 8'h00;
Ins_Reg[241] = 8'h0f;
Ins_Reg[242] = 8'h0f;
Ins_Reg[243] = 8'h13;
Ins_Reg[244] = 8'h00;
Ins_Reg[245] = 8'h85;
Ins_Reg[246] = 8'h2f;
Ins_Reg[247] = 8'h03;
Ins_Reg[248] = 8'h00;
Ins_Reg[249] = 8'h0f;
Ins_Reg[250] = 8'h0f;
Ins_Reg[251] = 8'h13;
Ins_Reg[252] = 8'h01;
Ins_Reg[253] = 8'h05;
Ins_Reg[254] = 8'h23;
Ins_Reg[255] = 8'h03;
Ins_Reg[256] = 8'h00;
Ins_Reg[257] = 8'h0f;
Ins_Reg[258] = 8'h0f;
Ins_Reg[259] = 8'h13;
Ins_Reg[260] = 8'h01;
Ins_Reg[261] = 8'h85;
Ins_Reg[262] = 8'h23;
Ins_Reg[263] = 8'h83;
    end
    always @(posedge clk or reset)
    begin
    if (reset)
        Instruction <= 0;
    else if (clk)
    begin
        if(!(IF_ID_write) && clk) begin
        Instruction[7:0] <= Instruction[7:0];
        Instruction[15:8] <= Instruction[15:8];
        Instruction[23:16] <= Instruction[23:16];
        Instruction[31:24] <= Instruction[31:24];
        end
        else begin
        Instruction[7:0] <= Ins_Reg[Instr_Address+ 2'b11];
        Instruction[15:8] <= Ins_Reg[Instr_Address + 2'b10];
        Instruction[23:16] <= Ins_Reg[Instr_Address + 1'b1];
        Instruction[31:24] <= Ins_Reg[Instr_Address];
        end
        end
    end    
    
endmodule